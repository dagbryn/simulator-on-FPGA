library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

package arith_lib is

  function log(x : std_logic_vector)
    return std_logic_vector;

  function exp(x : std_logic_vector)
    return std_logic_vector;

  function sin(x : std_logic_vector)
    return std_logic_vector;

  function add(a, b : std_logic_vector)
    return std_logic_vector;

  function to_float(a, pos : signed)
    return std_logic_vector;

  function to_fixed(a : std_logic_vector; size, pos : unsigned)
    return signed;

  function multiply(a, b : std_logic_vector)
    return std_logic_vector;

end package arith_lib;

package body arith_lib is

  function log(x : std_logic_vector)
    return std_logic_vector is
    type rom_type is array(0 to 23) of unsigned(23 downto 0);
    variable rom : rom_type := (
      -- log(10) log(1.1) log(1.01)
      x"B17218", x"67CC8F", x"391FEF", x"1E2707",
      x"0F8518", x"07E0A6", x"03F815", x"01FE02",
      x"00FF80", x"007FE0", x"003FF8", x"001FFE",
      x"000FFF", x"0007FF", x"0003FF", x"0001FF",
      x"0000FF", x"00007F", x"00003F", x"00001F",
      x"00000F", x"000007", x"000003", x"000001"
      );
    variable tmp           : signed(31 downto 0) := (others => '0');
    variable result        : std_logic_vector(31 downto 0);
    variable mant, mant_in : unsigned(24 downto 0);
    variable mant_out      : unsigned(24 downto 0);
    variable expn          : signed(7 downto 0);
    variable pos           : signed(7 downto 0);
    variable mant20 : signed(22 downto 0);
  begin
    mant_in  := "01" & unsigned(x(22 downto 0));
    mant_out := '0' & rom(0);
    expn     := signed(x(30 downto 23)) - 127;
    for j in 1 to 23 loop
      mant := mant_in + shift_right(mant_in, j);
      if mant(mant'high) = '0' then
        mant_in  := mant;
        mant_out := mant_out - rom(j);
      end if;
    end loop;
    --if expn > 0 then
    tmp := expn * ('0' & signed(rom(0)(23 downto 1)));
    tmp := (tmp(tmp'high-1 downto 0) & '0') + ('0' & signed(mant_out));
    pos    := x"07";
    mant20 := tmp(tmp'high downto tmp'high-22);
    result := to_float(mant20, pos);
  return result;
end;

function exp(x : std_logic_vector)
  return std_logic_vector is
  type rom_type is array(0 to 1023) of std_logic_vector(31 downto 0);
  variable rom_low : rom_type := (
    x"3F800000", x"3F800120", x"3F800240", x"3F800360",
    x"3F800480", x"3F8005A0", x"3F8006C0", x"3F8007E0",
    x"3F800900", x"3F800A20", x"3F800B40", x"3F800C61",
    x"3F800D81", x"3F800EA1", x"3F800FC1", x"3F8010E1",
    x"3F801201", x"3F801321", x"3F801442", x"3F801562",
    x"3F801682", x"3F8017A2", x"3F8018C2", x"3F8019E3",
    x"3F801B03", x"3F801C23", x"3F801D43", x"3F801E64",
    x"3F801F84", x"3F8020A4", x"3F8021C4", x"3F8022E5",
    x"3F802405", x"3F802525", x"3F802646", x"3F802766",
    x"3F802886", x"3F8029A7", x"3F802AC7", x"3F802BE8",
    x"3F802D08", x"3F802E28", x"3F802F49", x"3F803069",
    x"3F80318A", x"3F8032AA", x"3F8033CA", x"3F8034EB",
    x"3F80360B", x"3F80372C", x"3F80384C", x"3F80396D",
    x"3F803A8D", x"3F803BAE", x"3F803CCE", x"3F803DEF",
    x"3F803F10", x"3F804030", x"3F804151", x"3F804271",
    x"3F804392", x"3F8044B2", x"3F8045D3", x"3F8046F4",
    x"3F804814", x"3F804935", x"3F804A56", x"3F804B76",
    x"3F804C97", x"3F804DB8", x"3F804ED8", x"3F804FF9",
    x"3F80511A", x"3F80523A", x"3F80535B", x"3F80547C",
    x"3F80559D", x"3F8056BD", x"3F8057DE", x"3F8058FF",
    x"3F805A20", x"3F805B40", x"3F805C61", x"3F805D82",
    x"3F805EA3", x"3F805FC4", x"3F8060E5", x"3F806205",
    x"3F806326", x"3F806447", x"3F806568", x"3F806689",
    x"3F8067AA", x"3F8068CB", x"3F8069EC", x"3F806B0D",
    x"3F806C2E", x"3F806D4F", x"3F806E70", x"3F806F91",
    x"3F8070B1", x"3F8071D2", x"3F8072F3", x"3F807415",
    x"3F807536", x"3F807657", x"3F807778", x"3F807899",
    x"3F8079BA", x"3F807ADB", x"3F807BFC", x"3F807D1D",
    x"3F807E3E", x"3F807F5F", x"3F808080", x"3F8081A1",
    x"3F8082C3", x"3F8083E4", x"3F808505", x"3F808626",
    x"3F808747", x"3F808868", x"3F80898A", x"3F808AAB",
    x"3F808BCC", x"3F808CED", x"3F808E0F", x"3F808F30",
    x"3F809051", x"3F809172", x"3F809294", x"3F8093B5",
    x"3F8094D6", x"3F8095F8", x"3F809719", x"3F80983A",
    x"3F80995C", x"3F809A7D", x"3F809B9E", x"3F809CC0",
    x"3F809DE1", x"3F809F02", x"3F80A024", x"3F80A145",
    x"3F80A267", x"3F80A388", x"3F80A4AA", x"3F80A5CB",
    x"3F80A6EC", x"3F80A80E", x"3F80A92F", x"3F80AA51",
    x"3F80AB72", x"3F80AC94", x"3F80ADB5", x"3F80AED7",
    x"3F80AFF9", x"3F80B11A", x"3F80B23C", x"3F80B35D",
    x"3F80B47F", x"3F80B5A0", x"3F80B6C2", x"3F80B7E4",
    x"3F80B905", x"3F80BA27", x"3F80BB48", x"3F80BC6A",
    x"3F80BD8C", x"3F80BEAD", x"3F80BFCF", x"3F80C0F1",
    x"3F80C213", x"3F80C334", x"3F80C456", x"3F80C578",
    x"3F80C699", x"3F80C7BB", x"3F80C8DD", x"3F80C9FF",
    x"3F80CB21", x"3F80CC42", x"3F80CD64", x"3F80CE86",
    x"3F80CFA8", x"3F80D0CA", x"3F80D1EB", x"3F80D30D",
    x"3F80D42F", x"3F80D551", x"3F80D673", x"3F80D795",
    x"3F80D8B7", x"3F80D9D9", x"3F80DAFA", x"3F80DC1C",
    x"3F80DD3E", x"3F80DE60", x"3F80DF82", x"3F80E0A4",
    x"3F80E1C6", x"3F80E2E8", x"3F80E40A", x"3F80E52C",
    x"3F80E64E", x"3F80E770", x"3F80E892", x"3F80E9B4",
    x"3F80EAD6", x"3F80EBF8", x"3F80ED1B", x"3F80EE3D",
    x"3F80EF5F", x"3F80F081", x"3F80F1A3", x"3F80F2C5",
    x"3F80F3E7", x"3F80F509", x"3F80F62C", x"3F80F74E",
    x"3F80F870", x"3F80F992", x"3F80FAB4", x"3F80FBD6",
    x"3F80FCF9", x"3F80FE1B", x"3F80FF3D", x"3F81005F",
    x"3F810182", x"3F8102A4", x"3F8103C6", x"3F8104E9",
    x"3F81060B", x"3F81072D", x"3F81084F", x"3F810972",
    x"3F810A94", x"3F810BB6", x"3F810CD9", x"3F810DFB",
    x"3F810F1E", x"3F811040", x"3F811162", x"3F811285",
    x"3F8113A7", x"3F8114CA", x"3F8115EC", x"3F81170E",
    x"3F811831", x"3F811953", x"3F811A76", x"3F811B98",
    x"3F811CBB", x"3F811DDD", x"3F811F00", x"3F812022",
    x"3F812145", x"3F812267", x"3F81238A", x"3F8124AD",
    x"3F8125CF", x"3F8126F2", x"3F812814", x"3F812937",
    x"3F812A5A", x"3F812B7C", x"3F812C9F", x"3F812DC2",
    x"3F812EE4", x"3F813007", x"3F81312A", x"3F81324C",
    x"3F81336F", x"3F813492", x"3F8135B4", x"3F8136D7",
    x"3F8137FA", x"3F81391D", x"3F813A3F", x"3F813B62",
    x"3F813C85", x"3F813DA8", x"3F813ECA", x"3F813FED",
    x"3F814110", x"3F814233", x"3F814356", x"3F814479",
    x"3F81459B", x"3F8146BE", x"3F8147E1", x"3F814904",
    x"3F814A27", x"3F814B4A", x"3F814C6D", x"3F814D90",
    x"3F814EB3", x"3F814FD6", x"3F8150F9", x"3F81521C",
    x"3F81533E", x"3F815461", x"3F815584", x"3F8156A7",
    x"3F8157CA", x"3F8158EE", x"3F815A11", x"3F815B34",
    x"3F815C57", x"3F815D7A", x"3F815E9D", x"3F815FC0",
    x"3F8160E3", x"3F816206", x"3F816329", x"3F81644C",
    x"3F81656F", x"3F816693", x"3F8167B6", x"3F8168D9",
    x"3F8169FC", x"3F816B1F", x"3F816C42", x"3F816D66",
    x"3F816E89", x"3F816FAC", x"3F8170CF", x"3F8171F3",
    x"3F817316", x"3F817439", x"3F81755C", x"3F817680",
    x"3F8177A3", x"3F8178C6", x"3F8179EA", x"3F817B0D",
    x"3F817C30", x"3F817D54", x"3F817E77", x"3F817F9A",
    x"3F8180BE", x"3F8181E1", x"3F818305", x"3F818428",
    x"3F81854B", x"3F81866F", x"3F818792", x"3F8188B6",
    x"3F8189D9", x"3F818AFD", x"3F818C20", x"3F818D44",
    x"3F818E67", x"3F818F8B", x"3F8190AE", x"3F8191D2",
    x"3F8192F5", x"3F819419", x"3F81953C", x"3F819660",
    x"3F819783", x"3F8198A7", x"3F8199CB", x"3F819AEE",
    x"3F819C12", x"3F819D35", x"3F819E59", x"3F819F7D",
    x"3F81A0A0", x"3F81A1C4", x"3F81A2E8", x"3F81A40B",
    x"3F81A52F", x"3F81A653", x"3F81A776", x"3F81A89A",
    x"3F81A9BE", x"3F81AAE2", x"3F81AC05", x"3F81AD29",
    x"3F81AE4D", x"3F81AF71", x"3F81B095", x"3F81B1B8",
    x"3F81B2DC", x"3F81B400", x"3F81B524", x"3F81B648",
    x"3F81B76C", x"3F81B88F", x"3F81B9B3", x"3F81BAD7",
    x"3F81BBFB", x"3F81BD1F", x"3F81BE43", x"3F81BF67",
    x"3F81C08B", x"3F81C1AF", x"3F81C2D3", x"3F81C3F7",
    x"3F81C51B", x"3F81C63F", x"3F81C763", x"3F81C887",
    x"3F81C9AB", x"3F81CACF", x"3F81CBF3", x"3F81CD17",
    x"3F81CE3B", x"3F81CF5F", x"3F81D083", x"3F81D1A7",
    x"3F81D2CB", x"3F81D3EF", x"3F81D513", x"3F81D638",
    x"3F81D75C", x"3F81D880", x"3F81D9A4", x"3F81DAC8",
    x"3F81DBEC", x"3F81DD10", x"3F81DE35", x"3F81DF59",
    x"3F81E07D", x"3F81E1A1", x"3F81E2C6", x"3F81E3EA",
    x"3F81E50E", x"3F81E632", x"3F81E757", x"3F81E87B",
    x"3F81E99F", x"3F81EAC4", x"3F81EBE8", x"3F81ED0C",
    x"3F81EE31", x"3F81EF55", x"3F81F079", x"3F81F19E",
    x"3F81F2C2", x"3F81F3E6", x"3F81F50B", x"3F81F62F",
    x"3F81F754", x"3F81F878", x"3F81F99C", x"3F81FAC1",
    x"3F81FBE5", x"3F81FD0A", x"3F81FE2E", x"3F81FF53",
    x"3F820077", x"3F82019C", x"3F8202C0", x"3F8203E5",
    x"3F820509", x"3F82062E", x"3F820752", x"3F820877",
    x"3F82099C", x"3F820AC0", x"3F820BE5", x"3F820D09",
    x"3F820E2E", x"3F820F53", x"3F821077", x"3F82119C",
    x"3F8212C1", x"3F8213E5", x"3F82150A", x"3F82162F",
    x"3F821753", x"3F821878", x"3F82199D", x"3F821AC2",
    x"3F821BE6", x"3F821D0B", x"3F821E30", x"3F821F55",
    x"3F822079", x"3F82219E", x"3F8222C3", x"3F8223E8",
    x"3F82250D", x"3F822631", x"3F822756", x"3F82287B",
    x"3F8229A0", x"3F822AC5", x"3F822BEA", x"3F822D0F",
    x"3F822E33", x"3F822F58", x"3F82307D", x"3F8231A2",
    x"3F8232C7", x"3F8233EC", x"3F823511", x"3F823636",
    x"3F82375B", x"3F823880", x"3F8239A5", x"3F823ACA",
    x"3F823BEF", x"3F823D14", x"3F823E39", x"3F823F5E",
    x"3F824083", x"3F8241A8", x"3F8242CD", x"3F8243F3",
    x"3F824518", x"3F82463D", x"3F824762", x"3F824887",
    x"3F8249AC", x"3F824AD1", x"3F824BF6", x"3F824D1C",
    x"3F824E41", x"3F824F66", x"3F82508B", x"3F8251B0",
    x"3F8252D6", x"3F8253FB", x"3F825520", x"3F825645",
    x"3F82576B", x"3F825890", x"3F8259B5", x"3F825ADA",
    x"3F825C00", x"3F825D25", x"3F825E4A", x"3F825F70",
    x"3F826095", x"3F8261BA", x"3F8262E0", x"3F826405",
    x"3F82652B", x"3F826650", x"3F826775", x"3F82689B",
    x"3F8269C0", x"3F826AE6", x"3F826C0B", x"3F826D31",
    x"3F826E56", x"3F826F7B", x"3F8270A1", x"3F8271C6",
    x"3F8272EC", x"3F827411", x"3F827537", x"3F82765D",
    x"3F827782", x"3F8278A8", x"3F8279CD", x"3F827AF3",
    x"3F827C18", x"3F827D3E", x"3F827E64", x"3F827F89",
    x"3F8280AF", x"3F8281D4", x"3F8282FA", x"3F828420",
    x"3F828545", x"3F82866B", x"3F828791", x"3F8288B6",
    x"3F8289DC", x"3F828B02", x"3F828C28", x"3F828D4D",
    x"3F828E73", x"3F828F99", x"3F8290BF", x"3F8291E4",
    x"3F82930A", x"3F829430", x"3F829556", x"3F82967C",
    x"3F8297A1", x"3F8298C7", x"3F8299ED", x"3F829B13",
    x"3F829C39", x"3F829D5F", x"3F829E85", x"3F829FAB",
    x"3F82A0D0", x"3F82A1F6", x"3F82A31C", x"3F82A442",
    x"3F82A568", x"3F82A68E", x"3F82A7B4", x"3F82A8DA",
    x"3F82AA00", x"3F82AB26", x"3F82AC4C", x"3F82AD72",
    x"3F82AE98", x"3F82AFBE", x"3F82B0E4", x"3F82B20A",
    x"3F82B330", x"3F82B456", x"3F82B57D", x"3F82B6A3",
    x"3F82B7C9", x"3F82B8EF", x"3F82BA15", x"3F82BB3B",
    x"3F82BC61", x"3F82BD87", x"3F82BEAE", x"3F82BFD4",
    x"3F82C0FA", x"3F82C220", x"3F82C346", x"3F82C46D",
    x"3F82C593", x"3F82C6B9", x"3F82C7DF", x"3F82C906",
    x"3F82CA2C", x"3F82CB52", x"3F82CC78", x"3F82CD9F",
    x"3F82CEC5", x"3F82CFEB", x"3F82D112", x"3F82D238",
    x"3F82D35E", x"3F82D485", x"3F82D5AB", x"3F82D6D2",
    x"3F82D7F8", x"3F82D91E", x"3F82DA45", x"3F82DB6B",
    x"3F82DC92", x"3F82DDB8", x"3F82DEDE", x"3F82E005",
    x"3F82E12B", x"3F82E252", x"3F82E378", x"3F82E49F",
    x"3F82E5C5", x"3F82E6EC", x"3F82E812", x"3F82E939",
    x"3F82EA60", x"3F82EB86", x"3F82ECAD", x"3F82EDD3",
    x"3F82EEFA", x"3F82F021", x"3F82F147", x"3F82F26E",
    x"3F82F394", x"3F82F4BB", x"3F82F5E2", x"3F82F708",
    x"3F82F82F", x"3F82F956", x"3F82FA7C", x"3F82FBA3",
    x"3F82FCCA", x"3F82FDF1", x"3F82FF17", x"3F83003E",
    x"3F830165", x"3F83028C", x"3F8303B2", x"3F8304D9",
    x"3F830600", x"3F830727", x"3F83084E", x"3F830974",
    x"3F830A9B", x"3F830BC2", x"3F830CE9", x"3F830E10",
    x"3F830F37", x"3F83105E", x"3F831184", x"3F8312AB",
    x"3F8313D2", x"3F8314F9", x"3F831620", x"3F831747",
    x"3F83186E", x"3F831995", x"3F831ABC", x"3F831BE3",
    x"3F831D0A", x"3F831E31", x"3F831F58", x"3F83207F",
    x"3F8321A6", x"3F8322CD", x"3F8323F4", x"3F83251B",
    x"3F832642", x"3F832769", x"3F832891", x"3F8329B8",
    x"3F832ADF", x"3F832C06", x"3F832D2D", x"3F832E54",
    x"3F832F7B", x"3F8330A3", x"3F8331CA", x"3F8332F1",
    x"3F833418", x"3F83353F", x"3F833667", x"3F83378E",
    x"3F8338B5", x"3F8339DC", x"3F833B04", x"3F833C2B",
    x"3F833D52", x"3F833E79", x"3F833FA1", x"3F8340C8",
    x"3F8341EF", x"3F834317", x"3F83443E", x"3F834565",
    x"3F83468D", x"3F8347B4", x"3F8348DC", x"3F834A03",
    x"3F834B2A", x"3F834C52", x"3F834D79", x"3F834EA1",
    x"3F834FC8", x"3F8350F0", x"3F835217", x"3F83533E",
    x"3F835466", x"3F83558D", x"3F8356B5", x"3F8357DC",
    x"3F835904", x"3F835A2C", x"3F835B53", x"3F835C7B",
    x"3F835DA2", x"3F835ECA", x"3F835FF1", x"3F836119",
    x"3F836241", x"3F836368", x"3F836490", x"3F8365B7",
    x"3F8366DF", x"3F836807", x"3F83692E", x"3F836A56",
    x"3F836B7E", x"3F836CA5", x"3F836DCD", x"3F836EF5",
    x"3F83701D", x"3F837144", x"3F83726C", x"3F837394",
    x"3F8374BC", x"3F8375E3", x"3F83770B", x"3F837833",
    x"3F83795B", x"3F837A83", x"3F837BAB", x"3F837CD2",
    x"3F837DFA", x"3F837F22", x"3F83804A", x"3F838172",
    x"3F83829A", x"3F8383C2", x"3F8384EA", x"3F838611",
    x"3F838739", x"3F838861", x"3F838989", x"3F838AB1",
    x"3F838BD9", x"3F838D01", x"3F838E29", x"3F838F51",
    x"3F839079", x"3F8391A1", x"3F8392C9", x"3F8393F1",
    x"3F839519", x"3F839641", x"3F83976A", x"3F839892",
    x"3F8399BA", x"3F839AE2", x"3F839C0A", x"3F839D32",
    x"3F839E5A", x"3F839F82", x"3F83A0AB", x"3F83A1D3",
    x"3F83A2FB", x"3F83A423", x"3F83A54B", x"3F83A673",
    x"3F83A79C", x"3F83A8C4", x"3F83A9EC", x"3F83AB14",
    x"3F83AC3D", x"3F83AD65", x"3F83AE8D", x"3F83AFB5",
    x"3F83B0DE", x"3F83B206", x"3F83B32E", x"3F83B457",
    x"3F83B57F", x"3F83B6A7", x"3F83B7D0", x"3F83B8F8",
    x"3F83BA21", x"3F83BB49", x"3F83BC71", x"3F83BD9A",
    x"3F83BEC2", x"3F83BFEB", x"3F83C113", x"3F83C23B",
    x"3F83C364", x"3F83C48C", x"3F83C5B5", x"3F83C6DD",
    x"3F83C806", x"3F83C92E", x"3F83CA57", x"3F83CB7F",
    x"3F83CCA8", x"3F83CDD1", x"3F83CEF9", x"3F83D022",
    x"3F83D14A", x"3F83D273", x"3F83D39B", x"3F83D4C4",
    x"3F83D5ED", x"3F83D715", x"3F83D83E", x"3F83D967",
    x"3F83DA8F", x"3F83DBB8", x"3F83DCE1", x"3F83DE09",
    x"3F83DF32", x"3F83E05B", x"3F83E184", x"3F83E2AC",
    x"3F83E3D5", x"3F83E4FE", x"3F83E627", x"3F83E74F",
    x"3F83E878", x"3F83E9A1", x"3F83EACA", x"3F83EBF3",
    x"3F83ED1B", x"3F83EE44", x"3F83EF6D", x"3F83F096",
    x"3F83F1BF", x"3F83F2E8", x"3F83F411", x"3F83F539",
    x"3F83F662", x"3F83F78B", x"3F83F8B4", x"3F83F9DD",
    x"3F83FB06", x"3F83FC2F", x"3F83FD58", x"3F83FE81",
    x"3F83FFAA", x"3F8400D3", x"3F8401FC", x"3F840325",
    x"3F84044E", x"3F840577", x"3F8406A0", x"3F8407C9",
    x"3F8408F2", x"3F840A1B", x"3F840B44", x"3F840C6E",
    x"3F840D97", x"3F840EC0", x"3F840FE9", x"3F841112",
    x"3F84123B", x"3F841364", x"3F84148E", x"3F8415B7",
    x"3F8416E0", x"3F841809", x"3F841932", x"3F841A5C",
    x"3F841B85", x"3F841CAE", x"3F841DD7", x"3F841F01",
    x"3F84202A", x"3F842153", x"3F84227D", x"3F8423A6",
    x"3F8424CF", x"3F8425F8", x"3F842722", x"3F84284B",
    x"3F842975", x"3F842A9E", x"3F842BC7", x"3F842CF1",
    x"3F842E1A", x"3F842F43", x"3F84306D", x"3F843196",
    x"3F8432C0", x"3F8433E9", x"3F843513", x"3F84363C",
    x"3F843766", x"3F84388F", x"3F8439B9", x"3F843AE2",
    x"3F843C0C", x"3F843D35", x"3F843E5F", x"3F843F88",
    x"3F8440B2", x"3F8441DB", x"3F844305", x"3F84442F",
    x"3F844558", x"3F844682", x"3F8447AB", x"3F8448D5",
    x"3F8449FF", x"3F844B28", x"3F844C52", x"3F844D7C",
    x"3F844EA5", x"3F844FCF", x"3F8450F9", x"3F845223",
    x"3F84534C", x"3F845476", x"3F8455A0", x"3F8456C9",
    x"3F8457F3", x"3F84591D", x"3F845A47", x"3F845B71",
    x"3F845C9A", x"3F845DC4", x"3F845EEE", x"3F846018",
    x"3F846142", x"3F84626C", x"3F846396", x"3F8464BF",
    x"3F8465E9", x"3F846713", x"3F84683D", x"3F846967",
    x"3F846A91", x"3F846BBB", x"3F846CE5", x"3F846E0F",
    x"3F846F39", x"3F847063", x"3F84718D", x"3F8472B7",
    x"3F8473E1", x"3F84750B", x"3F847635", x"3F84775F",
    x"3F847889", x"3F8479B3", x"3F847ADD", x"3F847C07",
    x"3F847D31", x"3F847E5B", x"3F847F85", x"3F8480B0",
    x"3F8481DA", x"3F848304", x"3F84842E", x"3F848558",
    x"3F848682", x"3F8487AD", x"3F8488D7", x"3F848A01",
    x"3F848B2B", x"3F848C55", x"3F848D80", x"3F848EAA",
    x"3F848FD4", x"3F8490FE", x"3F849229", x"3F849353"
    );
  variable rom_high : rom_type := (
    x"3282D314", x"32878171", x"328C5AAF", x"32916057",
    x"329693FF", x"329BF74E", x"32A18BF7", x"32A753BE",
    x"32AD5079", x"32B3840B", x"32B9F06C", x"32C097A3",
    x"32C77BCC", x"32CE9F15", x"32D603C0", x"32DDAC24",
    x"32E59AAD", x"32EDD1DE", x"32F65450", x"32FF24B5",
    x"330422EC", x"3308DD4D", x"330DC2FD", x"3312D589",
    x"3318168C", x"331D87AF", x"33232AAC", x"3329014A",
    x"332F0D63", x"333550E1", x"333BCDBF", x"3342860B",
    x"33497BE5", x"3350B180", x"33582926", x"335FE532",
    x"3367E818", x"33703460", x"3378CCAB", x"3380D9D8",
    x"33857621", x"338A3CA5", x"338F2EE8", x"33944E79",
    x"33999CF9", x"339F1C15", x"33A4CD8A", x"33AAB325",
    x"33B0CEC4", x"33B72256", x"33BDAFDC", x"33C47968",
    x"33CB8120", x"33D2C93D", x"33DA540E", x"33E223F6",
    x"33EA3B6C", x"33F29D02", x"33FB4B5D", x"3402249E",
    x"3406CCBD", x"340B9F84", x"34109E79", x"3415CB31",
    x"341B2751", x"3420B488", x"3426749B", x"342C6959",
    x"343294A7", x"3438F876", x"343F96CF", x"344671C7",
    x"344D8B8B", x"3454E65A", x"345C8487", x"3464687D",
    x"346C94B9", x"34750BD2", x"347DD076", x"348372B6",
    x"348826C9", x"348D05F1", x"349211BA", x"34974BBB",
    x"349CB59C", x"34A25115", x"34A81FEA", x"34AE23F3",
    x"34B45F16", x"34BAD34D", x"34C182A3", x"34C86F35",
    x"34CF9B33", x"34D708E3", x"34DEBA9F", x"34E6B2D6",
    x"34EEF40D", x"34F780E2", x"35002E04", x"3504C427",
    x"3509844D", x"350E6FF7", x"351388B3", x"3518D01F",
    x"351E47E7", x"3523F1C4", x"3529CF82", x"352FE2FC",
    x"35362E1F", x"353CB2E7", x"35437366", x"354A71BE",
    x"3551B025", x"355930E8", x"3560F664", x"35690310",
    x"35715978", x"3579FC40", x"35817711", x"358618FA",
    x"358AE552", x"358FDD9E", x"35950370", x"359A5869",
    x"359FDE39", x"35A596A1", x"35AB836E", x"35B1A681",
    x"35B801CC", x"35BE9750", x"35C56924", x"35CC7970",
    x"35D3CA70", x"35DB5E75", x"35E337E5", x"35EB593B",
    x"35F3C50A", x"35FC7DFD", x"3602C36B", x"36077138",
    x"360C49E1", x"36114EEF", x"361681F8", x"361BE4A1",
    x"3621789F", x"36273FB6", x"362D3BB9", x"36336E8D",
    x"3639DA29", x"36408095", x"364763EA", x"364E8659",
    x"3655EA21", x"365D919A", x"36657F30", x"366DB565",
    x"367636D3", x"367F062A", x"3684131A", x"3688CCEA",
    x"368DB204", x"3692C3F5", x"36980457", x"369D74D3",
    x"36A31723", x"36A8ED0E", x"36AEF86E", x"36B53B2C",
    x"36BBB744", x"36C26EC1", x"36C963C6", x"36D09884",
    x"36D80F45", x"36DFCA64", x"36E7CC55", x"36F0179E",
    x"36F8AEE2", x"3700CA6B", x"37056627", x"370A2C18",
    x"370F1DC3", x"37143CB8", x"37198A95", x"371F0908",
    x"3724B9CF", x"372A9EB5", x"3730B999", x"37370C6A",
    x"373D9927", x"374461E2", x"374B68C3", x"3752B001",
    x"375A39EB", x"376208E3", x"376A1F62", x"37727FF6",
    x"377B2D47", x"3782150A", x"3786BC9A", x"378B8ECC",
    x"37908D29", x"3795B943", x"379B14BD", x"37A0A14B",
    x"37A660AD", x"37AC54B5", x"37B27F45", x"37B8E251",
    x"37BF7FDF", x"37C65A05", x"37CD72EF", x"37D4CCDD",
    x"37DC6A21", x"37E44D24", x"37EC7866", x"37F4EE7C",
    x"37FDB213", x"380362F9", x"3808167C", x"380CF50F",
    x"3812003D", x"3817399E", x"381CA2D9", x"38223DA6",
    x"38280BC9", x"382E0F19", x"3834497E", x"383ABCEF",
    x"38416B78", x"38485736", x"384F8258", x"3856EF25",
    x"385E9FF5", x"38669737", x"386ED772", x"38776340",
    x"38801EAB", x"3884B442", x"388973D6", x"388E5EE9",
    x"3893770A", x"3898BDD4", x"389E34F3", x"38A3DE23",
    x"38A9BB2E", x"38AFCDED", x"38B6184F", x"38BC9C50",
    x"38C35C00", x"38CA5981", x"38D1970B", x"38D916E7",
    x"38E0DB75", x"38E8E72B", x"38F13C93", x"38F9DE52",
    x"39016791", x"390608EC", x"390AD4B1", x"390FCC64",
    x"3914F199", x"391A45EE", x"391FCB16", x"392582CE",
    x"392B6EE5", x"3931913D", x"3937EBC4", x"393E807F",
    x"39455182", x"394C60F5", x"3953B115", x"395B4432",
    x"39631CB1", x"396B3D0E", x"3973A7DB", x"397C5FC3",
    x"3982B3C3", x"39876101", x"398C3916", x"39913D8A",
    x"39966FF3", x"399BD1F8", x"39A1654B", x"39A72BB0",
    x"39AD26FC", x"39B35912", x"39B9C3E9", x"39C06989",
    x"39C74C0C", x"39CE6D9F", x"39D5D085", x"39DD7713",
    x"39E563B6", x"39ED98F0", x"39F61959", x"39FEE7A2",
    x"3A04034A", x"3A08BC89", x"3A0DA10D", x"3A12B263",
    x"3A17F224", x"3A1D61F9", x"3A23039D", x"3A28D8D5",
    x"3A2EE37C", x"3A35257A", x"3A3BA0CA", x"3A42577A",
    x"3A494BA9", x"3A507F8B", x"3A57F567", x"3A5FAF9A",
    x"3A67B094", x"3A6FFAE0", x"3A78911C", x"3A80BB00",
    x"3A85562E", x"3A8A1B8E", x"3A8F0CA1", x"3A942AF9",
    x"3A997833", x"3A9EF5FE", x"3AA4A616", x"3AAA8A48",
    x"3AB0A471", x"3AB6F680", x"3ABD8274", x"3AC44A60",
    x"3ACB5069", x"3AD296C8", x"3ADA1FCB", x"3AE1EDD3",
    x"3AEA035A", x"3AF262EE", x"3AFB0F35", x"3B020577",
    x"3B06AC78", x"3B0B7E17", x"3B107BDA", x"3B15A756",
    x"3B1B022C", x"3B208E10", x"3B264CC2", x"3B2C4014",
    x"3B3269E7", x"3B38CC2F", x"3B3F68F2", x"3B464246",
    x"3B4D5A57", x"3B54B363", x"3B5C4FBE", x"3B6431CF",
    x"3B6C5C17", x"3B74D129", x"3B7D93B4", x"3B83533E",
    x"3B880631", x"3B8CE42F", x"3B91EEC2", x"3B972783",
    x"3B9C9019", x"3BA22A39", x"3BA7F7AB", x"3BADFA43",
    x"3BB433E9", x"3BBAA694", x"3BC15450", x"3BC83F39",
    x"3BCF6980", x"3BD6D569", x"3BDE854E", x"3BE67B9C",
    x"3BEEBAD9", x"3BF745A2", x"3C000F55", x"3C04A45F",
    x"3C096361", x"3C0E4DDE", x"3C136562", x"3C18AB8B",
    x"3C1E2203", x"3C23CA85", x"3C29A6DC", x"3C2FB8E1",
    x"3C360282", x"3C3C85BB", x"3C43449C", x"3C4A4148",
    x"3C517DF3", x"3C58FCEA", x"3C60C08A", x"3C68CB49",
    x"3C711FB2", x"3C79C068", x"3C815813", x"3C85F8E0",
    x"3C8AC412", x"3C8FBB2D", x"3C94DFC4", x"3C9A3376",
    x"3C9FB7F4", x"3CA56EFD", x"3CAB5A5F", x"3CB17BFA",
    x"3CB7D5BF", x"3CBE69B0", x"3CC539E2", x"3CCC487E",
    x"3CD397BD", x"3CDB29F2", x"3CE30180", x"3CEB20E4",
    x"3CF38AB0", x"3CFC418C", x"3D02A41D", x"3D0750CC",
    x"3D0C284C", x"3D112C26", x"3D165DF1", x"3D1BBF50",
    x"3D2151F8", x"3D2717AD", x"3D2D1241", x"3D334399",
    x"3D39ADAC", x"3D405280", x"3D47342F", x"3D4E54E8",
    x"3D55B6EC", x"3D5D5C90", x"3D654840", x"3D6D7C7E",
    x"3D75FBE2", x"3D7EC91D", x"3D83F37C", x"3D88AC2B",
    x"3D8D9019", x"3D92A0D3", x"3D97DFF3", x"3D9D4F22",
    x"3DA2F019", x"3DA8C49E", x"3DAECE8C", x"3DB50FCA",
    x"3DBB8A54", x"3DC24036", x"3DC93390", x"3DD06695",
    x"3DD7DB8C", x"3DDF94D2", x"3DE794D7", x"3DEFDE25",
    x"3DF8735A", x"3E00AB97", x"3E054638", x"3E0A0B05",
    x"3E0EFB81", x"3E14193C", x"3E1965D4", x"3E1EE2F6",
    x"3E249260", x"3E2A75DD", x"3E308F4B", x"3E36E098",
    x"3E3D6BC4", x"3E4432E0", x"3E4B3812", x"3E527D92",
    x"3E5A05AE", x"3E61D2C7", x"3E69E756", x"3E7245E9",
    x"3E7AF126", x"3E81F5E6", x"3E869C59", x"3E8B6D64",
    x"3E906A8E", x"3E95956B", x"3E9AEF9E", x"3EA07AD7",
    x"3EA638D9", x"3EAC2B74", x"3EB2548B", x"3EB8B60F",
    x"3EBF5207", x"3EC62A8A", x"3ECD41C1", x"3ED499EC",
    x"3EDC355D", x"3EE4167E", x"3EEC3FCB", x"3EF4B3DA",
    x"3EFD7558", x"3F034385", x"3F07F5E8", x"3F0CD351",
    x"3F11DD4A", x"3F17156A", x"3F1C7D5A", x"3F2216CF",
    x"3F27E38F", x"3F2DE56F", x"3F341E56", x"3F3A903C",
    x"3F413D2B", x"3F482740", x"3F4F50AC", x"3F56BBB1",
    x"3F5E6AAA", x"3F666004", x"3F6E9E45", x"3F772808",
    x"3F800000", x"3F84947D", x"3F8952EF", x"3F8E3CD4",
    x"3F9353BD", x"3F989944", x"3F9E0F14", x"3FA3B6E9",
    x"3FA9928C", x"3FAFA3D8", x"3FB5ECB8", x"3FBC6F29",
    x"3FC32D3C", x"3FCA2911", x"3FD164DF", x"3FD8E2EF",
    x"3FE0A5A2", x"3FE8AF6A", x"3FF102D4", x"3FF9A282",
    x"40014897", x"4005E8D6", x"400AB375", x"400FA9F8",
    x"4014CDF1", x"401A2100", x"401FA4D5", x"40255B2F",
    x"402B45DC", x"403166BB", x"4037BFBD", x"403E52E5",
    x"40452246", x"404C3009", x"40537E68", x"405B0FB5",
    x"4062E653", x"406B04BE", x"40736D87", x"407C2359",
    x"40829479", x"40874099", x"408C1785", x"40911AC5",
    x"40964BF0", x"409BACAB", x"40A13EA8", x"40A703AC",
    x"40ACFD89", x"40B32E23", x"40B99771", x"40C03B79",
    x"40C71C56", x"40CE3C35", x"40D59D56", x"40DD420F",
    x"40E52CCD", x"40ED600F", x"40F5DE6F", x"40FEAA9D",
    x"4103E3B0", x"41089BCE", x"410D7F26", x"41128F45",
    x"4117CDC4", x"411D3C4D", x"4122DC97", x"4128B06A",
    x"412EB99E", x"4134FA1D", x"413B73E0", x"414228F5",
    x"41491B7A", x"41504DA2", x"4157C1B5", x"415F7A0E",
    x"4167791E", x"416FC16D", x"4178559B", x"41809C2F",
    x"41853643", x"4189FA7E", x"418EEA63", x"41940781",
    x"41995376", x"419ECFF1", x"41A47EAC", x"41AA6175",
    x"41B07A28", x"41B6CAB3", x"41BD5516", x"41C41B63",
    x"41CB1FBD", x"41D2645F", x"41D9EB94", x"41E1B7BE",
    x"41E9CB55", x"41F228E8", x"41FAD31B", x"4201E657",
    x"42068C3B", x"420B5CB3", x"42105944", x"42158383",
    x"421ADD11", x"422067A1", x"422624F3", x"422C16D8",
    x"42323F31", x"42389FF2", x"423F3B20", x"424612D0",
    x"424D292E", x"42548078", x"425C1B00", x"4263FB2F",
    x"426C2382", x"4274968E", x"427D5700", x"428333CE",
    x"4287E5A1", x"428CC275", x"4291CBD3", x"42970354",
    x"429C6A9E", x"42A20368", x"42A7CF75", x"42ADD09D",
    x"42B408C5", x"42BA79E6", x"42C12609", x"42C80F4A",
    x"42CF37DA", x"42D6A1FC", x"42DE5009", x"42E64470",
    x"42EE81B4", x"42F70A71", x"42FFE15A", x"4304849E",
    x"4309427E", x"430E2BCD", x"43134219", x"431886FF",
    x"431DFC28", x"4323A34F", x"43297E3F", x"432F8ED1",
    x"4335D6F0", x"433C589A", x"434315DE", x"434A10DD",
    x"43514BCD", x"4358C8F8", x"43608ABD", x"4368938F",
    x"4370E5F9", x"4379849F", x"4381391D", x"4385D8CE",
    x"438AA2DA", x"438F98C5", x"4394BC20", x"439A0E8D",
    x"439F91B9", x"43A54763", x"43AB315A", x"43B1517E",
    x"43B7A9BE", x"43BE3C1B", x"43C50AAC", x"43CC1797",
    x"43D36516", x"43DAF57B", x"43E2CB29", x"43EAE89B",
    x"43F35063", x"43FC0529", x"440284D7", x"44073068",
    x"440C06BF", x"44110966", x"441639F2", x"441B9A07",
    x"44212B5A", x"4426EFAD", x"442CE8D3", x"443318B0",
    x"44398139", x"44402476", x"44470480", x"444E2384",
    x"445583C3", x"445D2792", x"4465115D", x"446D43A4",
    x"4475C100", x"447E8C1F", x"4483D3E6", x"44888B73",
    x"448D6E36", x"44927DB9", x"4497BB98", x"449D297A",
    x"44A2C917", x"44A89C38", x"44AEA4B3", x"44B4E472",
    x"44BB5D6F", x"44C211B6", x"44C90366", x"44D034B2",
    x"44D7A7E0", x"44DF5F4C", x"44E75D68", x"44EFA4B9",
    x"44F837E0", x"45008CC9", x"45052650", x"4509E9F9",
    x"450ED947", x"4513F5C8", x"4519411B", x"451EBCED",
    x"45246AFB", x"452A4D0F", x"45306507", x"4536B4D1",
    x"453D3E6B", x"454403E8", x"454B076C", x"45524B2F",
    x"4559D17D", x"45619CB8", x"4569AF58", x"45720BEA",
    x"457AB514", x"4581D6CA", x"45867C20", x"458B4C04",
    x"459047FC", x"4595719C", x"459ACA87", x"45A0546D",
    x"45A6110F", x"45AC023D", x"45B229DA", x"45B889D8",
    x"45BF243B", x"45C5FB19", x"45CD109E", x"45D46707",
    x"45DC00A7", x"45E3DFE4", x"45EC073D", x"45F47946",
    x"45FD38AC", x"46032419", x"4607D55C", x"460CB19B",
    x"4611BA5F", x"4616F140", x"461C57E4", x"4621F002",
    x"4627BB5E", x"462DBBCE", x"4633F338", x"463A6393",
    x"46410EE9", x"4647F756", x"464F1F0B", x"4656884A",
    x"465E356C", x"466628DE", x"466E6526", x"4676ECDD",
    x"467FC2B8", x"468474C1", x"4689320F", x"468E1AC8",
    x"46933078", x"469874BC", x"469DE93E", x"46A38FB8",
    x"46A969F4", x"46AF79CC", x"46B5C12B", x"46BC420E",
    x"46C2FE83", x"46C9F8AC", x"46D132BF", x"46D8AF04",
    x"46E06FDB", x"46E877B7", x"46F0C922", x"46F966C0",
    x"470129A4", x"4705C8C8", x"470A9241", x"470F8794",
    x"4714AA52", x"4719FC1B", x"471F7E9E", x"47253399",
    x"472B1CDC", x"47313C43", x"473793C1", x"473E2555",
    x"4744F315", x"474BFF28", x"47534BC8", x"475ADB44",
    x"4762B002", x"476ACC7C", x"47733342", x"477BE6FD",
    x"47827537", x"47872038", x"478BF5FB", x"4790F809",
    x"479627F6", x"479B8767", x"47A1180F", x"47A6DBB1",
    x"47ACD41F", x"47B3033F", x"47B96B04", x"47C00D75",
    x"47C6ECAC", x"47CE0AD6", x"47D56A33", x"47DD0D18",
    x"47E4F5F0", x"47ED273C", x"47F5A394", x"47FE6DA6",
    x"4803C41E", x"48087B1A", x"480D5D47", x"48126C2F",
    x"4817A96D", x"481D16A9", x"4822B59A", x"48288808",
    x"482E8FCB", x"4834CECA", x"483B4701", x"4841FA7A",
    x"4848EB55", x"48501BC5", x"48578E0F", x"485F448E",
    x"486741B5", x"486F8809", x"48781A29", x"48807D66",
    x"4885165F", x"4889D977", x"488EC82D", x"4893E411",
    x"48992EC2", x"489EA9EC", x"48A4574C", x"48AA38AC",
    x"48B04FE9", x"48B69EF1", x"48BD27C4", x"48C3EC71",
    x"48CAEF1D", x"48D23201", x"48D9B769", x"48E181B6",
    x"48E9935E", x"48F1EEF0", x"48FA9710", x"4901C73E",
    x"49066C06", x"490B3B56", x"491036B6", x"49155FB8",
    x"491AB7FF", x"4920413B", x"4925FD2D", x"492BEDA6",
    x"49321486", x"493873C0", x"493F0D59", x"4945E366",
    x"494CF812", x"49544D9A", x"495BE650", x"4963C49C",
    x"496BEAFB", x"49745C01", x"497D1A5B", x"49831466",
    x"4987C519", x"498CA0C3", x"4991A8EC", x"4996DF2E",
    x"499C452D", x"49A1DC9F", x"49A7A74A", x"49ADA701",
    x"49B3DDAD", x"49BA4D42", x"49C0F7CC", x"49C7DF66",
    x"49CF063F", x"49D66E9B", x"49DE1AD1", x"49E60D50",
    x"49EE489B", x"49F6CF4D", x"49FFA419", x"4A0464E5",
    x"4A0921A2", x"4A0E09C5", x"4A131ED9", x"4A18627B",
    x"4A1DD656", x"4A237C23", x"4A2955AC", x"4A2F64CA",
    x"4A35AB69", x"4A3C2B84", x"4A42E72B", x"4A49E07E",
    x"4A5119B3", x"4A589513", x"4A6054FC", x"4A685BE2",
    x"4A70AC4F", x"4A7948E4", x"4A811A2E", x"4A85B8C4",
    x"4A8A81AA", x"4A8F7665", x"4A949886", x"4A99E9AC",
    x"4A9F6B86", x"4AA51FD2", x"4AAB085F", x"4AB1270B",
    x"4AB77DC6", x"4ABE0E92", x"4AC4DB81", x"4ACBE6BB",
    x"4AD3327C", x"4ADAC111", x"4AE294DE", x"4AEAB05F",
    x"4AF31624", x"4AFBC8D5", x"4B026599", x"4B07100B",
    x"4B0BE53A", x"4B10E6AE", x"4B1615FC", x"4B1B74C8",
    x"4B2104C5", x"4B26C7B7", x"4B2CBF6F", x"4B32EDD0",
    x"4B3954D1", x"4B3FF677", x"4B46D4DC", x"4B4DF22B",
    x"4B5550A6", x"4B5CF2A1", x"4B64DA87", x"4B6D0AD8",
    x"4B75862B", x"4B7E4F30", x"4B83B457", x"4B886AC3",
    x"4B8D4C5A", x"4B925AA8", x"4B979745", x"4B9D03DB",
    x"4BA2A21F", x"4BA873DB", x"4BAE7AE5", x"4BB4B925",
    x"4BBB3095", x"4BC1E341", x"4BC8D348", x"4BD002DB",
    x"4BD77440", x"4BDF29D4", x"4BE72605", x"4BEF6B5C",
    x"4BF7FC75", x"4C006E04", x"4C050671", x"4C09C8F6",
    x"4C0EB715", x"4C13D25D", x"4C191C6C", x"4C1E96EE",
    x"4C24439F", x"4C2A244B", x"4C303ACE", x"4C368914",
    x"4C3D111E", x"4C43D4FC", x"4C4AD6D2", x"4C5218D7",
    x"4C599D58", x"4C6166B6", x"4C697767", x"4C71D1F9"
    );
  variable xh, xl : integer range 0 to 1023;
begin
  xl := to_integer(unsigned(x(x'low+9 downto x'low)));
  xh := to_integer(unsigned(x(19 downto 10)));
  return multiply(rom_high(xh),
                  rom_low(xl));
end;

function sin(x : std_logic_vector)
  return std_logic_vector is
  type rom_type is array(0 to 1023) of std_logic_vector(31 downto 0);
  variable rom : rom_type := (
    x"00000000", x"00646EC8", x"00C8DD82", x"012D4C1C",
    x"0191BA88", x"01F628B6", x"025A9696", x"02BF0419",
    x"03237131", x"0387DDCC", x"03EC49DC", x"0450B550",
    x"04B5201B", x"05198A2C", x"057DF373", x"05E25BE2",
    x"0646C368", x"06AB29F7", x"070F8F7E", x"0773F3EE",
    x"07D85739", x"083CB94D", x"08A11A1C", x"09057997",
    x"0969D7AE", x"09CE3451", x"0A328F70", x"0A96E8FE",
    x"0AFB40E9", x"0B5F9722", x"0BC3EB9B", x"0C283E43",
    x"0C8C8F0B", x"0CF0DDE4", x"0D552ABE", x"0DB9758A",
    x"0E1DBE37", x"0E8204B8", x"0EE648FB", x"0F4A8AF3",
    x"0FAECA8F", x"101307BF", x"10774275", x"10DB7AA1",
    x"113FB034", x"11A3E31E", x"1208134F", x"126C40B8",
    x"12D06B4A", x"133492F5", x"1398B7AB", x"13FCD95A",
    x"1460F7F4", x"14C5136A", x"15292BAC", x"158D40AA",
    x"15F15256", x"1655609F", x"16B96B77", x"171D72CE",
    x"17817694", x"17E576BA", x"18497330", x"18AD6BE8",
    x"191160D2", x"197551DE", x"19D93EFD", x"1A3D281F",
    x"1AA10D36", x"1B04EE31", x"1B68CB02", x"1BCCA399",
    x"1C3077E6", x"1C9447DA", x"1CF81366", x"1D5BDA7A",
    x"1DBF9D07", x"1E235AFE", x"1E87144F", x"1EEAC8EB",
    x"1F4E78C3", x"1FB223C6", x"2015C9E6", x"20796B13",
    x"20DD073F", x"21409E59", x"21A43052", x"2207BD1B",
    x"226B44A5", x"22CEC6E0", x"233243BC", x"2395BB2C",
    x"23F92D1E", x"245C9984", x"24C0004F", x"2523616F",
    x"2586BCD4", x"25EA1271", x"264D6234", x"26B0AC0F",
    x"2713EFF3", x"27772DD0", x"27DA6598", x"283D9739",
    x"28A0C2A6", x"2903E7D0", x"296706A6", x"29CA1F19",
    x"2A2D311B", x"2A903C9C", x"2AF3418C", x"2B563FDD",
    x"2BB9377E", x"2C1C2862", x"2C7F1278", x"2CE1F5B2",
    x"2D44D200", x"2DA7A753", x"2E0A759B", x"2E6D3CC9",
    x"2ECFFCCF", x"2F32B59D", x"2F956723", x"2FF81153",
    x"305AB41D", x"30BD4F72", x"311FE343", x"31826F81",
    x"31E4F41C", x"32477106", x"32A9E62E", x"330C5386",
    x"336EB8FF", x"33D1168A", x"34336C17", x"3495B997",
    x"34F7FEFB", x"355A3C34", x"35BC7132", x"361E9DE8",
    x"3680C245", x"36E2DE3A", x"3744F1B8", x"37A6FCB0",
    x"3808FF13", x"386AF8D2", x"38CCE9DE", x"392ED227",
    x"3990B19F", x"39F28837", x"3A5455DE", x"3AB61A87",
    x"3B17D622", x"3B7988A0", x"3BDB31F2", x"3C3CD20A",
    x"3C9E68D7", x"3CFFF64A", x"3D617A56", x"3DC2F4EB",
    x"3E2465F9", x"3E85CD72", x"3EE72B47", x"3F487F68",
    x"3FA9C9C7", x"400B0A55", x"406C4102", x"40CD6DC0",
    x"412E9080", x"418FA933", x"41F0B7C9", x"4251BC34",
    x"42B2B665", x"4313A64D", x"43748BDD", x"43D56705",
    x"443637B8", x"4496FDE6", x"44F7B980", x"45586A77",
    x"45B910BD", x"4619AC42", x"467A3CF7", x"46DAC2CE",
    x"473B3DB8", x"479BADA6", x"47FC1289", x"485C6C52",
    x"48BCBAF3", x"491CFE5C", x"497D367E", x"49DD634B",
    x"4A3D84B5", x"4A9D9AAB", x"4AFDA520", x"4B5DA404",
    x"4BBD9748", x"4C1D7EDF", x"4C7D5AB9", x"4CDD2AC7",
    x"4D3CEEFA", x"4D9CA745", x"4DFC5397", x"4E5BF3E3",
    x"4EBB8819", x"4F1B102A", x"4F7A8C09", x"4FD9FBA7",
    x"50395EF3", x"5098B5E1", x"50F80061", x"51573E64",
    x"51B66FDC", x"521594BA", x"5274ACF0", x"52D3B86F",
    x"5332B727", x"5391A90B", x"53F08E0C", x"544F661B",
    x"54AE312A", x"550CEF29", x"556BA00B", x"55CA43C1",
    x"5628DA3C", x"5687636D", x"56E5DF46", x"57444DB9",
    x"57A2AEB7", x"58010231", x"585F4818", x"58BD805F",
    x"591BAAF7", x"5979C7D0", x"59D7D6DE", x"5A35D810",
    x"5A93CB59", x"5AF1B0AA", x"5B4F87F5", x"5BAD512B",
    x"5C0B0C3E", x"5C68B91F", x"5CC657C0", x"5D23E813",
    x"5D816A08", x"5DDEDD92", x"5E3C42A2", x"5E99992A",
    x"5EF6E11B", x"5F541A67", x"5FB144FF", x"600E60D6",
    x"606B6DDD", x"60C86C05", x"61255B41", x"61823B81",
    x"61DF0CB8", x"623BCED7", x"629881CF", x"62F52594",
    x"6351BA15", x"63AE3F46", x"640AB518", x"64671B7C",
    x"64C37264", x"651FB9C2", x"657BF188", x"65D819A8",
    x"66343213", x"66903ABB", x"66EC3392", x"67481C8A",
    x"67A3F595", x"67FFBEA4", x"685B77A9", x"68B72096",
    x"6912B95E", x"696E41F1", x"69C9BA42", x"6A252243",
    x"6A8079E5", x"6ADBC11B", x"6B36F7D6", x"6B921E08",
    x"6BED33A4", x"6C48389B", x"6CA32CDF", x"6CFE1063",
    x"6D58E317", x"6DB3A4EF", x"6E0E55DB", x"6E68F5CF",
    x"6EC384BC", x"6F1E0295", x"6F786F4A", x"6FD2CACF",
    x"702D1516", x"70874E0F", x"70E175AF", x"713B8BE6",
    x"719590A7", x"71EF83E3", x"7249658E", x"72A33599",
    x"72FCF3F6", x"7356A097", x"73B03B6F", x"7409C470",
    x"74633B8C", x"74BCA0B5", x"7515F3DE", x"756F34F8",
    x"75C863F6", x"762180CA", x"767A8B67", x"76D383BE",
    x"772C69C2", x"77853D66", x"77DDFE9B", x"7836AD53",
    x"788F4982", x"78E7D31A", x"79404A0C", x"7998AE4B",
    x"79F0FFCA", x"7A493E7B", x"7AA16A51", x"7AF9833D",
    x"7B518932", x"7BA97C23", x"7C015C01", x"7C5928C1",
    x"7CB0E253", x"7D0888AA", x"7D601BBA", x"7DB79B74",
    x"7E0F07CB", x"7E6660B1", x"7EBDA619", x"7F14D7F5",
    x"7F6BF639", x"7FC300D6", x"8019F7BF", x"8070DAE7",
    x"80C7AA41", x"811E65BE", x"81750D52", x"81CBA0F0",
    x"82222089", x"82788C10", x"82CEE379", x"832526B6",
    x"837B55B9", x"83D17076", x"842776DF", x"847D68E6",
    x"84D3467F", x"85290F9D", x"857EC431", x"85D4642F",
    x"8629EF8A", x"867F6634", x"86D4C820", x"872A1542",
    x"877F4D8B", x"87D470F0", x"88297F61", x"887E78D4",
    x"88D35D3A", x"89282C86", x"897CE6AB", x"89D18B9D",
    x"8A261B4E", x"8A7A95B1", x"8ACEFAB9", x"8B234A59",
    x"8B778484", x"8BCBA92D", x"8C1FB847", x"8C73B1C5",
    x"8CC7959B", x"8D1B63BB", x"8D6F1C18", x"8DC2BEA5",
    x"8E164B56", x"8E69C21E", x"8EBD22F0", x"8F106DBE",
    x"8F63A27C", x"8FB6C11E", x"9009C996", x"905CBBD8",
    x"90AF97D6", x"91025D84", x"91550CD6", x"91A7A5BE",
    x"91FA2830", x"924C941F", x"929EE97F", x"92F12842",
    x"9343505C", x"939561C0", x"93E75C62", x"94394035",
    x"948B0D2C", x"94DCC33B", x"952E6256", x"957FEA6E",
    x"95D15B79", x"9622B569", x"9673F832", x"96C523C8",
    x"9716381D", x"97673526", x"97B81AD5", x"9808E91F",
    x"98599FF7", x"98AA3F50", x"98FAC71E", x"994B3755",
    x"999B8FE8", x"99EBD0CB", x"9A3BF9F1", x"9A8C0B4E",
    x"9ADC04D6", x"9B2BE67D", x"9B7BB035", x"9BCB61F4",
    x"9C1AFBAB", x"9C6A7D50", x"9CB9E6D6", x"9D093831",
    x"9D587154", x"9DA79234", x"9DF69AC3", x"9E458AF6",
    x"9E9462C1", x"9EE32218", x"9F31C8EE", x"9F805737",
    x"9FCECCE7", x"A01D29F2", x"A06B6E4D", x"A0B999EA",
    x"A107ACBE", x"A155A6BD", x"A1A387DA", x"A1F1500A",
    x"A23EFF41", x"A28C9573", x"A2DA1294", x"A3277698",
    x"A374C172", x"A3C1F318", x"A40F0B7C", x"A45C0A94",
    x"A4A8F053", x"A4F5BCAE", x"A5426F98", x"A58F0906",
    x"A5DB88EC", x"A627EF3F", x"A6743BF1", x"A6C06EF9",
    x"A70C8849", x"A75887D7", x"A7A46D96", x"A7F0397A",
    x"A83BEB79", x"A8878386", x"A8D30196", x"A91E659D",
    x"A969AF8F", x"A9B4DF62", x"A9FFF508", x"AA4AF077",
    x"AA95D1A4", x"AAE09882", x"AB2B4506", x"AB75D724",
    x"ABC04ED1", x"AC0AAC02", x"AC54EEAC", x"AC9F16C1",
    x"ACE92438", x"AD331705", x"AD7CEF1C", x"ADC6AC72",
    x"AE104EFB", x"AE59D6AD", x"AEA3437C", x"AEEC955C",
    x"AF35CC42", x"AF7EE824", x"AFC7E8F5", x"B010CEAB",
    x"B059993A", x"B0A24897", x"B0EADCB6", x"B133558D",
    x"B17BB311", x"B1C3F536", x"B20C1BF1", x"B2542737",
    x"B29C16FD", x"B2E3EB37", x"B32BA3DC", x"B37340DF",
    x"B3BAC235", x"B40227D4", x"B44971B1", x"B4909FC0",
    x"B4D7B1F7", x"B51EA84A", x"B56582AF", x"B5AC411B",
    x"B5F2E383", x"B63969DB", x"B67FD41A", x"B6C62234",
    x"B70C541E", x"B75269CE", x"B7986339", x"B7DE4053",
    x"B8240113", x"B869A56D", x"B8AF2D57", x"B8F498C6",
    x"B939E7AF", x"B97F1A07", x"B9C42FC5", x"BA0928DC",
    x"BA4E0544", x"BA92C4F0", x"BAD767D7", x"BB1BEDED",
    x"BB605729", x"BBA4A37F", x"BBE8D2E6", x"BC2CE552",
    x"BC70DAB9", x"BCB4B311", x"BCF86E4F", x"BD3C0C69",
    x"BD7F8D55", x"BDC2F107", x"BE063775", x"BE496096",
    x"BE8C6C5F", x"BECF5AC5", x"BF122BBE", x"BF54DF40",
    x"BF977540", x"BFD9EDB5", x"C01C4894", x"C05E85D3",
    x"C0A0A567", x"C0E2A746", x"C1248B67", x"C16651BF",
    x"C1A7FA43", x"C1E984EB", x"C22AF1AB", x"C26C4079",
    x"C2AD714D", x"C2EE841A", x"C32F78D8", x"C3704F7C",
    x"C3B107FD", x"C3F1A250", x"C4321E6C", x"C4727C46",
    x"C4B2BBD5", x"C4F2DD0E", x"C532DFE8", x"C572C459",
    x"C5B28A57", x"C5F231D9", x"C631BAD3", x"C671253E",
    x"C6B0710E", x"C6EF9E3A", x"C72EACB9", x"C76D9C80",
    x"C7AC6D86", x"C7EB1FC1", x"C829B328", x"C86827B0",
    x"C8A67D51", x"C8E4B401", x"C922CBB5", x"C960C466",
    x"C99E9E07", x"C9DC5892", x"CA19F3FB", x"CA57703A",
    x"CA94CD44", x"CAD20B11", x"CB0F2997", x"CB4C28CC",
    x"CB8908A8", x"CBC5C920", x"CC026A2C", x"CC3EEBC1",
    x"CC7B4DD8", x"CCB79066", x"CCF3B362", x"CD2FB6C2",
    x"CD6B9A7F", x"CDA75E8D", x"CDE302E5", x"CE1E877D",
    x"CE59EC4B", x"CE953147", x"CED05667", x"CF0B5BA3",
    x"CF4640F1", x"CF810648", x"CFBBAB9F", x"CFF630ED",
    x"D030962A", x"D06ADB4B", x"D0A50048", x"D0DF0518",
    x"D118E9B2", x"D152AE0E", x"D18C5222", x"D1C5D5E5",
    x"D1FF394E", x"D2387C56", x"D2719EF2", x"D2AAA11A",
    x"D2E382C5", x"D31C43EB", x"D354E483", x"D38D6483",
    x"D3C5C3E4", x"D3FE029C", x"D43620A3", x"D46E1DF1",
    x"D4A5FA7C", x"D4DDB63C", x"D5155128", x"D54CCB38",
    x"D5842464", x"D5BB5CA2", x"D5F273EA", x"D6296A34",
    x"D6603F77", x"D696F3AB", x"D6CD86C8", x"D703F8C4",
    x"D73A4998", x"D770793B", x"D7A687A5", x"D7DC74CD",
    x"D81240AB", x"D847EB38", x"D87D746A", x"D8B2DC39",
    x"D8E8229D", x"D91D478E", x"D9524B04", x"D9872CF6",
    x"D9BBED5D", x"D9F08C2F", x"DA250966", x"DA5964F9",
    x"DA8D9EE0", x"DAC1B713", x"DAF5AD89", x"DB29823C",
    x"DB5D3522", x"DB90C634", x"DBC4356A", x"DBF782BC",
    x"DC2AAE22", x"DC5DB794", x"DC909F0A", x"DCC3647D",
    x"DCF607E4", x"DD288939", x"DD5AE872", x"DD8D2589",
    x"DDBF4075", x"DDF1392E", x"DE230FAE", x"DE54C3ED",
    x"DE8655E2", x"DEB7C586", x"DEE912D1", x"DF1A3DBD",
    x"DF4B4640", x"DF7C2C55", x"DFACEFF2", x"DFDD9111",
    x"E00E0FAB", x"E03E6BB7", x"E06EA52E", x"E09EBC09",
    x"E0CEB040", x"E0FE81CD", x"E12E30A6", x"E15DBCC7",
    x"E18D2626", x"E1BC6CBC", x"E1EB9083", x"E21A9173",
    x"E2496F85", x"E2782AB1", x"E2A6C2F1", x"E2D5383D",
    x"E3038A8D", x"E331B9DC", x"E35FC621", x"E38DAF56",
    x"E3BB7574", x"E3E91873", x"E416984D", x"E443F4F9",
    x"E4712E73", x"E49E44B2", x"E4CB37AF", x"E4F80764",
    x"E524B3CA", x"E5513CD9", x"E57DA28B", x"E5A9E4DA",
    x"E5D603BD", x"E601FF30", x"E62DD729", x"E6598BA4",
    x"E6851C99", x"E6B08A01", x"E6DBD3D6", x"E706FA11",
    x"E731FCAB", x"E75CDB9F", x"E78796E4", x"E7B22E75",
    x"E7DCA24B", x"E806F260", x"E8311EAC", x"E85B272A",
    x"E8850BD3", x"E8AECCA0", x"E8D8698B", x"E901E28E",
    x"E92B37A2", x"E95468C1", x"E97D75E5", x"E9A65F07",
    x"E9CF2420", x"E9F7C52C", x"EA204222", x"EA489AFE",
    x"EA70CFB8", x"EA98E04B", x"EAC0CCB1", x"EAE894E3",
    x"EB1038DB", x"EB37B893", x"EB5F1405", x"EB864B2B",
    x"EBAD5DFF", x"EBD44C7B", x"EBFB1699", x"EC21BC52",
    x"EC483DA1", x"EC6E9A81", x"EC94D2EA", x"ECBAE6D8",
    x"ECE0D643", x"ED06A128", x"ED2C477E", x"ED51C942",
    x"ED77266D", x"ED9C5EF8", x"EDC172E0", x"EDE6621D",
    x"EE0B2CAA", x"EE2FD282", x"EE54539E", x"EE78AFF9",
    x"EE9CE78E", x"EEC0FA57", x"EEE4E84F", x"EF08B16F",
    x"EF2C55B3", x"EF4FD514", x"EF732F8E", x"EF96651A",
    x"EFB975B4", x"EFDC6156", x"EFFF27FB", x"F021C99D",
    x"F0444637", x"F0669DC4", x"F088D03E", x"F0AADDA0",
    x"F0CCC5E5", x"F0EE8908", x"F1102703", x"F1319FD1",
    x"F152F36D", x"F17421D2", x"F1952AFB", x"F1B60EE3",
    x"F1D6CD84", x"F1F766DA", x"F217DAE0", x"F2382990",
    x"F25852E5", x"F27856DB", x"F298356D", x"F2B7EE96",
    x"F2D78250", x"F2F6F097", x"F3163967", x"F3355CBA",
    x"F3545A8B", x"F37332D6", x"F391E596", x"F3B072C7",
    x"F3CEDA63", x"F3ED1C65", x"F40B38CA", x"F4292F8D",
    x"F44700A8", x"F464AC18", x"F48231D7", x"F49F91E2",
    x"F4BCCC33", x"F4D9E0C6", x"F4F6CF98", x"F51398A2",
    x"F5303BE1", x"F54CB950", x"F56910EC", x"F58542AF",
    x"F5A14E95", x"F5BD349A", x"F5D8F4BA", x"F5F48EF0",
    x"F6100338", x"F62B518E", x"F64679EE", x"F6617C53",
    x"F67C58B9", x"F6970F1C", x"F6B19F79", x"F6CC09CA",
    x"F6E64E0D", x"F7006C3C", x"F71A6453", x"F7343650",
    x"F74DE22D", x"F76767E8", x"F780C77B", x"F79A00E3",
    x"F7B3141C", x"F7CC0122", x"F7E4C7F2", x"F7FD6887",
    x"F815E2DE", x"F82E36F3", x"F84664C2", x"F85E6C48",
    x"F8764D81", x"F88E0868", x"F8A59CFB", x"F8BD0B36",
    x"F8D45315", x"F8EB7495", x"F9026FB2", x"F9194468",
    x"F92FF2B4", x"F9467A93", x"F95CDC01", x"F97316FA",
    x"F9892B7B", x"F99F1981", x"F9B4E109", x"F9CA820E",
    x"F9DFFC8E", x"F9F55086", x"FA0A7DF1", x"FA1F84CE",
    x"FA346517", x"FA491ECB", x"FA5DB1E7", x"FA721E66",
    x"FA866446", x"FA9A8384", x"FAAE7C1C", x"FAC24E0B",
    x"FAD5F950", x"FAE97DE5", x"FAFCDBC9", x"FB1012F8",
    x"FB232370", x"FB360D2D", x"FB48D02D", x"FB5B6C6D",
    x"FB6DE1E9", x"FB8030A0", x"FB92588D", x"FBA459AF",
    x"FBB63402", x"FBC7E785", x"FBD97433", x"FBEADA0B",
    x"FBFC1909", x"FC0D312C", x"FC1E226F", x"FC2EECD2",
    x"FC3F9051", x"FC500CE9", x"FC606299", x"FC70915D",
    x"FC809933", x"FC907A19", x"FCA0340C", x"FCAFC70A",
    x"FCBF3310", x"FCCE781C", x"FCDD962C", x"FCEC8D3D",
    x"FCFB5D4D", x"FD0A0659", x"FD188860", x"FD26E35F",
    x"FD351755", x"FD43243D", x"FD510A18", x"FD5EC8E2",
    x"FD6C6099", x"FD79D13C", x"FD871AC8", x"FD943D3A",
    x"FDA13892", x"FDAE0CCE", x"FDBAB9EA", x"FDC73FE5",
    x"FDD39EBE", x"FDDFD672", x"FDEBE6FF", x"FDF7D064",
    x"FE03929F", x"FE0F2DAD", x"FE1AA18E", x"FE25EE3F",
    x"FE3113BF", x"FE3C120C", x"FE46E924", x"FE519905",
    x"FE5C21AE", x"FE66831E", x"FE70BD52", x"FE7AD04A",
    x"FE84BC03", x"FE8E807C", x"FE981DB3", x"FEA193A8",
    x"FEAAE258", x"FEB409C2", x"FEBD09E5", x"FEC5E2BF",
    x"FECE944F", x"FED71E94", x"FEDF818C", x"FEE7BD37",
    x"FEEFD192", x"FEF7BE9C", x"FEFF8455", x"FF0722BB",
    x"FF0E99CC", x"FF15E989", x"FF1D11EF", x"FF2412FD",
    x"FF2AECB3", x"FF319F10", x"FF382A12", x"FF3E8DB8",
    x"FF44CA01", x"FF4ADEED", x"FF50CC7A", x"FF5692A8",
    x"FF5C3176", x"FF61A8E2", x"FF66F8EC", x"FF6C2194",
    x"FF7122D8", x"FF75FCB7", x"FF7AAF31", x"FF7F3A45",
    x"FF839DF3", x"FF87DA39", x"FF8BEF17", x"FF8FDC8D",
    x"FF93A29A", x"FF97413C", x"FF9AB875", x"FF9E0843",
    x"FFA130A5", x"FFA4319B", x"FFA70B25", x"FFA9BD43",
    x"FFAC47F3", x"FFAEAB36", x"FFB0E70A", x"FFB2FB71",
    x"FFB4E868", x"FFB6ADF1", x"FFB84C0B", x"FFB9C2B5",
    x"FFBB11F0", x"FFBC39BB", x"FFBD3A16", x"FFBE1301",
    x"FFBEC47B", x"FFBF4E85", x"FFBFB11E", x"FFBFEC47"
    );
begin
  return ('0' & rom(to_integer(unsigned(x(x'low+9 downto x'low) xor (x'low+9 downto x'low => x(x'high-1)))))(31 downto 1))
    xor (31 downto 0 => x(x'high));
-- return ('0' & rom(to_integer(unsigned(x(9 downto 0) xor (9 downto 0 =>x(10)))))(31 downto 1))
--   xor (31 downto 0 => x(11));
end;

function add(a, b : std_logic_vector)
  return std_logic_vector is
  variable m_a, m_b, tmp_m : unsigned(24 downto 0);
  variable e_a, e_b, tmp_e : unsigned(8 downto 0);
  variable s_a, s_b, tmp_s : std_logic;
  variable i               : natural;
begin
  s_a := a(31); s_b := b(31);
  e_a := '0' & unsigned(a(30 downto 23)); e_b := '0' & unsigned(b(30 downto 23));
  m_a := "01" & unsigned(a(22 downto 0)); m_b := "01" & unsigned(b(22 downto 0));
  if e_a < e_b or (e_a = e_b and m_a < m_b) then  -- swap a,b
    s_a := b(31); s_b := a(31);
    e_a := '0' & unsigned(b(30 downto 23)); e_b := '0' & unsigned(a(30 downto 23));
    m_a := "01" & unsigned(b(22 downto 0)); m_b := "01" & unsigned(a(22 downto 0));
  end if;

  m_b := shift_right(m_b, to_integer(e_a - e_b));

  if s_a = s_b then
    m_a := m_a + m_b;
  else
    m_a := m_a - m_b;
  end if;
-- end of arg b

  e_a := e_a + 1;
  for j in 1 to 5 loop
    i := 2**(5-j);
    if m_a(m_a'high downto m_a'high-i+1) = (m_a'high downto m_a'high-i+1 => '0') then
      m_a := shift_left(m_a, i);
      e_a := e_a - i;
    end if;
  end loop;
  return s_a & std_logic_vector(e_a(7 downto 0)) & std_logic_vector(m_a(23 downto 1));
end;

function to_float(a, pos : signed)
  return std_logic_vector is
  variable m    : signed(a'high-a'low downto 0);
  variable expn : signed(pos'high-pos'low downto 0);
  variable i    : natural;
--  variable result : std_logic_vector(31 downto 0);
begin
  m    := abs(a);
  expn := pos;
  for j in 1 to 5 loop
    i := 2**(5-j);
    if m(m'high downto m'high-i+1) = (m'high downto m'high-i+1 => '0') then
      m    := shift_left(m, i);
      expn := expn - i;
    end if;
  end loop;
  return a(a'high) & std_logic_vector(expn+127) &
    std_logic_vector(m(m'high-1 downto 0)) & (22-m'high downto 0 => '0');
end;

function to_fixed(a : std_logic_vector; size, pos : unsigned)
  return signed is
  variable mant : signed(24 downto 0);
  variable expn : signed(7 downto 0);
  variable sign : std_logic;
begin
  sign := a(a'high);
  expn := signed(a(a'high-1 downto a'high-8));
  mant := signed("01" & a(22 downto 0));
  if signed(pos)-expn > -125 then
    mant := shift_right(mant, to_integer(signed(pos)-expn+125));
  end if;
  if sign = '1' then
    mant := -mant;
  end if;
  return mant(24 downto 5);             --to_integer(size));
end;

function multiply (a, b : std_logic_vector)
  return std_logic_vector is
  variable tmp  : unsigned(41 downto 0) := (others => '0');
  variable mant : unsigned(24 downto 0);
  variable expn : signed(8 downto 0);
begin
  tmp  := unsigned('1' & a(22 downto 0)) * unsigned('1' & b(22 downto 6));
  mant := tmp(tmp'high downto tmp'high-24);

  expn := signed('0' & a(30 downto 23)) + signed('0' & b(30 downto 23)) - 127;
  if mant(mant'high) = '1' then
    mant := '0' & tmp(tmp'high downto tmp'high-23);
    expn := expn + 1;
  end if;
  if expn(8) = '1' then
    expn := (others => '0');
  end if;

  return (a(31) xor b(31)) & std_logic_vector(expn(7 downto 0)) & std_logic_vector(mant(22 downto 0));
end;

end package body arith_lib;
